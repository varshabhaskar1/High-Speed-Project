module CLA_24bmod(a,b,sum,c_0);

input [24:0]a,b;

input c_0;

output [24:0]sum;

//output c_6;

wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,g0,g1,g2,g3,g4,g5,g6,g7,g8,g9,g10,g11,g12,g13,g14,g15,g16,g17,g18,g19,g20,g21,g22,g23,g24;

wire c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24;

assign

p0=a[0]^b[0],

p1=a[1]^b[1],

p2=a[2]^b[2],

p3=a[3]^b[3],

p4=a[4]^b[4],

p5=a[5]^b[5],

p6=a[6]^b[6],

p7=a[7]^b[7],

p8=a[8]^b[8],

p9=a[9]^b[9],

p10=a[10]^b[10],

p11=a[11]^b[11],

p12=a[12]^b[12],

p13=a[13]^b[13],

p14=a[14]^b[14],

p15=a[15]^b[15],


p16=a[16]^b[16],

p17=a[17]^b[17],

p18=a[18]^b[18],

p19=a[19]^b[19],

p20=a[20]^b[20],

p21=a[21]^b[21],

p22=a[22]^b[22],

p23=a[23]^b[23],
p24=a[24]^b[24],


g0=a[0]&b[0],

g1=a[1]&b[1],

g2=a[2]&b[2],

g3=a[3]&b[3],

g4=a[4]&b[4],

g5=a[5]&b[5],
g6=a[6]&b[6],

g7=a[7]&b[7],

g8=a[8]&b[8],

g9=a[9]&b[9],

g10=a[10]&b[10],

g11=a[11]&b[11],
g12=a[12]&b[12],

g13=a[13]&b[13],

g14=a[14]&b[14],

g15=a[15]&b[15],
g16=a[16]&b[16],

g17=a[17]&b[17],

g18=a[18]&b[18],

g19=a[19]&b[19],

g20=a[20]&b[20],

g21=a[21]&b[21],
g22=a[22]&b[22],

g23=a[23]&b[23];

g24=a[24]&b[24];

assign

c1=g0|(p0&c_0),

c2=g1|(p1&g0)|(p1&p0&c_0),

c3=g2|(p2&g1)|(p2&p1&g0)|(p2&p1&p0&c_0),

c4=g3|(p3&g2)|(p3&p2&g1)|(p3&p2&p1&g0)|(p3&p2&p1&p0&c_0),

c5=g4|(p4&g3)|(p4&p3&g2)|(p4&p3&p2&g1)|(p4&p3&p2&p1&g0)|(p4&p3&p2&p1&p0&c_0),
c6=g5|(p5&g4)|(p5&p4&g3)|( p5&p4&p3&g2 ) | ( p5&p4&p3&p2&g1) | (p5&p4&p3&p2&p1&g0) | (p5&p4&p3&p2&p1&p0&c_0),
c7= g6|(p6&g5)|(p6&p5&g4)|(p6&p5&p4&g3) | (p6&p5&p4&p3&g2) | (p6&p5&p4&p3&p2&g1) | (p6&p5&p4&p3&p2&p1&g0) | (p6&p5&p4&p3&p2&p1&p0&c_0 ),
c8=g7|(p7&g6) | (p7&p6&g5) |(p7 & p6 & p5 & g4) | (p7&p6&p5&p4&g3) | (p7&p6&p5&p4&p3&g2) | (p7&p6&p5&p4&p3&p2&g1) | (p7&p6&p5&p4&p3&p2&p1&g0) | (p7&p6&p5&p4&p3&p2&p1&p0&c_0 ),
c9=g8|(p8&g7)|(p8&p7&g6)|(p8&p7&p6&g5)|(p8&p7&p6&p5&g4)|(p8&p7&p6&p5&p4&g3)|(p8&p7&p6&p5&p4&p3&g2)|(p8&p7&p6&p5&p4&p3&p2&g1)|(p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p8&p7&p6&p5&p4&p3&p2&p1&p0&c_0),
c10=g9|(p9&g8)|(p9&p8&g7)|(p9&p8&p7&g6)|(p9&p8&p7&p6&g5)|(p9&p8&p7&p6&p5&g4)|(p9&p8&p7&p6&p5&p4&g3)|(p9&p8&p7&p6&p5&p4&p3&g2)|(p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c11=g10|p10&g9|(p10&p9&g8)|(p10&p9&p8&g7)|(p10&p9&p8&p7&g6)|(p10&p9&p8&p7&p6&g5)|(p10&p9&p8&p7&p6&p5&g4)|(p10&p9&p8&p7&p6&p5&p4&g3)|(p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c12=g11|p11&g10|p11&p10&g9|(p11&p10&p9&g8)|(p11&p10&p9&p8&g7)|(p11&p10&p9&p8&p7&g6)|(p11&p10&p9&p8&p7&p6&g5)|(p11&p10&p9&p8&p7&p6&p5&g4)|(p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c13=g12|p12&g11|p12&p11&g10|p12&p11&p10&g9|(p12&p11&p10&p9&g8)|(p12&p11&p10&p9&p8&g7)|(p12&p11&p10&p9&p8&p7&g6)|(p12&p11&p10&p9&p8&p7&p6&g5)|(p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c14=g13|(p13&g12)|(p13&p12&g11)|(p13&p12&p11&g10)|(p13&p12&p11&p10&g9)|(p13&p12&p11&p10&p9&g8)|(p13&p12&p11&p10&p9&p8&g7)|(p13&p12&p11&p10&p9&p8&p7&g6)|(p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c15=g14|(p14&g13)|(p14&p13&g12)|(p14&p13&p12&g11)|(p14&p13&p12&p11&g10)|(p14&p13&p12&p11&p10&g9)|(p14&p13&p12&p11&p10&p9&g8)|(p14&p13&p12&p11&p10&p9&p8&g7)|(p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c16=g15|(p15&g14)|(p15&p14&g13)|(p15&p14&p13&g12)|(p15&p14&p13&p12&g11)|(p15&p14&p13&p12&p11&g10)|(p15&p14&p13&p12&p11&p10&g9)|(p15&p14&p13&p12&p11&p10&p9&g8)|(p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c17=g16|(p16&g15)|(p16&p15&g14)|(p16&p15&p14&g13)|(p16&p15&p14&p13&g12)|(p16&p15&p14&p13&p12&g11)|(p16&p15&p14&p13&p12&p11&g10)|(p16&p15&p14&p13&p12&p11&p10&g9)|(p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c18=g17|(p17&p16&g15)|(p17&p16&p15&g14)|(p17&p16&p15&p14&g13)|(p17&p16&p15&p14&p13&g12)|(p17&p16&p15&p14&p13&p12&g11)|(p17&p16&p15&p14&p13&p12&p11&g10)|(p17&p16&p15&p14&p13&p12&p11&p10&g9)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c19=g18|(p18&g17)|(p18&p17&p16&g15)|(p18&p17&p16&p15&g14)|(p18&p17&p16&p15&p14&g13)|(p18&p17&p16&p15&p14&p13&g12)|(p18&p17&p16&p15&p14&p13&p12&g11)|(p18&p17&p16&p15&p14&p13&p12&p11&g10)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&g9)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c20=g19|(p19&g18)|(p19&p18&g17)|(p19&p18&p17&p16&g15)|(p19&p18&p17&p16&p15&g14)|(p19&p18&p17&p16&p15&p14&g13)|(p19&p18&p17&p16&p15&p14&p13&g12)|(p19&p18&p17&p16&p15&p14&p13&p12&g11)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&g10)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&g9)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),
c21=g20|(p20&g19)|(p20&p19&g18)|(p20&p19&p18&g17)|(p20&p19&p18&p17&p16&g15)|(p20&p19&p18&p17&p16&p15&g14)|(p20&p19&p18&p17&p16&p15&p14&g13)|(p20&p19&p18&p17&p16&p15&p14&p13&g12)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&g11)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&g10)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&g9)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),


c22=g21|(p21&g20)|(p21&p20&g19)|(p21&p20&p19&g18)|(p21&p20&p19&p18&g17)|(p21&p20&p19&p18&p17&p16&g15)|(p21&p20&p19&p18&p17&p16&p15&g14)|(p21&p20&p19&p18&p17&p16&p15&p14&g13)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&g12)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&g11)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&g10)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&g9)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),

c23=g22|(p22&g21)|(p22&p21&g20)|(p22&p21&p20&g19)|(p22&p21&p20&p19&g18)|(p22&p21&p20&p19&p18&g17)|(p22&p21&p20&p19&p18&p17&p16&g15)|(p22&p21&p20&p19&p18&p17&p16&p15&g14)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&g13)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&g12)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&g11)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&g10)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&g9)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0),

c24=g23|(p23&g22)|(p23&p22&g21)|(p23&p22&p21&g20)|(p23&p22&p21&p20&g19)|(p22&p21&p20&p19&g18)|(p23&p22&p21&p20&p19&p18&g17)|(p23&p22&p21&p20&p19&p18&p17&p16&g15)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&g14)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&g13)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&g12)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&g11)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&g10)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&g9)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&g8)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&g7)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&g6)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&g5)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&g4)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&g3)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&g2)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&g1)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&g0)|(p23&p22&p21&p20&p19&p18&p17&p16&p15&p14&p13&p12&p11&p10&p9&p8&p7&p6&p5&p4&p3&p2&p1&c_0);







assign

sum[0]=p0^c_0,

sum[1]=p1^c1,

sum[2]=p2^c2,

sum[3]=p3^c3,

sum[4]=p4^c4,

sum[5]=p5^c5,
sum[6]=p6^c6,
sum[7]=p7^c7,

sum[8]=p8^c8,

sum[9]=p9^c9,

sum[10]=p10^c10,

sum[11]=p11^c11,
sum[12]=p12^c12,

sum[13]=p13^c13,

sum[14]=p4^c14,

sum[15]=p15^c15,
sum[16]=p16^c16,
sum[17]=p17^c17,

sum[18]=p18^c18,

sum[19]=p19^c19,

sum[20]=p20^c20,

sum[21]=p21^c21,
sum[22]=p22^c22,

sum[23]=p23^c23;
sum[24]=p24^c24;

//c_6=c6;

endmodule




